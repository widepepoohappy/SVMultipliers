`timescale 10ns/1ns
module ANDoperator (input wire [7:0] A, 
 [7:0] B,
                  output wire [63:0] Out);
assign Out[0] = A[0] & B[0];
assign Out[1] = A[1] & B[0];
assign Out[2] = A[2] & B[0];
assign Out[3] = A[3] & B[0];
assign Out[4] = A[4] & B[0];
assign Out[5] = A[5] & B[0];
assign Out[6] = A[6] & B[0];
assign Out[7] = A[7] & B[0];
assign Out[8] = A[0] & B[1];
assign Out[9] = A[1] & B[1];
assign Out[10] = A[2] & B[1];
assign Out[11] = A[3] & B[1];
assign Out[12] = A[4] & B[1];
assign Out[13] = A[5] & B[1];
assign Out[14] = A[6] & B[1];
assign Out[15] = A[7] & B[1];
assign Out[16] = A[0] & B[2];
assign Out[17] = A[1] & B[2];
assign Out[18] = A[2] & B[2];
assign Out[19] = A[3] & B[2];
assign Out[20] = A[4] & B[2];
assign Out[21] = A[5] & B[2];
assign Out[22] = A[6] & B[2];
assign Out[23] = A[7] & B[2];
assign Out[24] = A[0] & B[3];
assign Out[25] = A[1] & B[3];
assign Out[26] = A[2] & B[3];
assign Out[27] = A[3] & B[3];
assign Out[28] = A[4] & B[3];
assign Out[29] = A[5] & B[3];
assign Out[30] = A[6] & B[3];
assign Out[31] = A[7] & B[3];
assign Out[32] = A[0] & B[4];
assign Out[33] = A[1] & B[4];
assign Out[34] = A[2] & B[4];
assign Out[35] = A[3] & B[4];
assign Out[36] = A[4] & B[4];
assign Out[37] = A[5] & B[4];
assign Out[38] = A[6] & B[4];
assign Out[39] = A[7] & B[4];
assign Out[40] = A[0] & B[5];
assign Out[41] = A[1] & B[5];
assign Out[42] = A[2] & B[5];
assign Out[43] = A[3] & B[5];
assign Out[44] = A[4] & B[5];
assign Out[45] = A[5] & B[5];
assign Out[46] = A[6] & B[5];
assign Out[47] = A[7] & B[5];
assign Out[48] = A[0] & B[6];
assign Out[49] = A[1] & B[6];
assign Out[50] = A[2] & B[6];
assign Out[51] = A[3] & B[6];
assign Out[52] = A[4] & B[6];
assign Out[53] = A[5] & B[6];
assign Out[54] = A[6] & B[6];
assign Out[55] = A[7] & B[6];
assign Out[56] = A[0] & B[7];
assign Out[57] = A[1] & B[7];
assign Out[58] = A[2] & B[7];
assign Out[59] = A[3] & B[7];
assign Out[60] = A[4] & B[7];
assign Out[61] = A[5] & B[7];
assign Out[62] = A[6] & B[7];
assign Out[63] = A[7] & B[7];
endmodule
