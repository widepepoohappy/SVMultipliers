`timescale 10ns/1ns
module Wallace_tree (input wire [64-1:0] INput,
                    (* keep *) output wire [16-1:0] WALLACEout [1:0]);


wire pp_s0_col0_row0;
wire pp_s0_col1_row0;
wire pp_s0_col1_row1;
wire pp_s0_col2_row0;
wire pp_s0_col2_row1;
wire pp_s0_col2_row2;
wire pp_s0_col3_row0;
wire pp_s0_col3_row1;
wire pp_s0_col3_row2;
wire pp_s0_col3_row3;
wire pp_s0_col4_row0;
wire pp_s0_col4_row1;
wire pp_s0_col4_row2;
wire pp_s0_col4_row3;
wire pp_s0_col4_row4;
wire pp_s0_col5_row0;
wire pp_s0_col5_row1;
wire pp_s0_col5_row2;
wire pp_s0_col5_row3;
wire pp_s0_col5_row4;
wire pp_s0_col5_row5;
wire pp_s0_col6_row0;
wire pp_s0_col6_row1;
wire pp_s0_col6_row2;
wire pp_s0_col6_row3;
wire pp_s0_col6_row4;
wire pp_s0_col6_row5;
wire pp_s0_col6_row6;
wire pp_s0_col7_row0;
wire pp_s0_col7_row1;
wire pp_s0_col7_row2;
wire pp_s0_col7_row3;
wire pp_s0_col7_row4;
wire pp_s0_col7_row5;
wire pp_s0_col7_row6;
wire pp_s0_col7_row7;
wire pp_s0_col8_row0;
wire pp_s0_col8_row1;
wire pp_s0_col8_row2;
wire pp_s0_col8_row3;
wire pp_s0_col8_row4;
wire pp_s0_col8_row5;
wire pp_s0_col8_row6;
wire pp_s0_col9_row0;
wire pp_s0_col9_row1;
wire pp_s0_col9_row2;
wire pp_s0_col9_row3;
wire pp_s0_col9_row4;
wire pp_s0_col9_row5;
wire pp_s0_col10_row0;
wire pp_s0_col10_row1;
wire pp_s0_col10_row2;
wire pp_s0_col10_row3;
wire pp_s0_col10_row4;
wire pp_s0_col11_row0;
wire pp_s0_col11_row1;
wire pp_s0_col11_row2;
wire pp_s0_col11_row3;
wire pp_s0_col12_row0;
wire pp_s0_col12_row1;
wire pp_s0_col12_row2;
wire pp_s0_col13_row0;
wire pp_s0_col13_row1;
wire pp_s0_col14_row0;

assign pp_s0_col0_row0 = INput[0];
assign pp_s0_col1_row0 = INput[1];
assign pp_s0_col1_row1 = INput[8];
assign pp_s0_col2_row0 = INput[2];
assign pp_s0_col2_row1 = INput[9];
assign pp_s0_col2_row2 = INput[16];
assign pp_s0_col3_row0 = INput[3];
assign pp_s0_col3_row1 = INput[10];
assign pp_s0_col3_row2 = INput[17];
assign pp_s0_col3_row3 = INput[24];
assign pp_s0_col4_row0 = INput[4];
assign pp_s0_col4_row1 = INput[11];
assign pp_s0_col4_row2 = INput[18];
assign pp_s0_col4_row3 = INput[25];
assign pp_s0_col4_row4 = INput[32];
assign pp_s0_col5_row0 = INput[5];
assign pp_s0_col5_row1 = INput[12];
assign pp_s0_col5_row2 = INput[19];
assign pp_s0_col5_row3 = INput[26];
assign pp_s0_col5_row4 = INput[33];
assign pp_s0_col5_row5 = INput[40];
assign pp_s0_col6_row0 = INput[6];
assign pp_s0_col6_row1 = INput[13];
assign pp_s0_col6_row2 = INput[20];
assign pp_s0_col6_row3 = INput[27];
assign pp_s0_col6_row4 = INput[34];
assign pp_s0_col6_row5 = INput[41];
assign pp_s0_col6_row6 = INput[48];
assign pp_s0_col7_row0 = INput[7];
assign pp_s0_col7_row1 = INput[14];
assign pp_s0_col7_row2 = INput[21];
assign pp_s0_col7_row3 = INput[28];
assign pp_s0_col7_row4 = INput[35];
assign pp_s0_col7_row5 = INput[42];
assign pp_s0_col7_row6 = INput[49];
assign pp_s0_col7_row7 = INput[56];
assign pp_s0_col8_row0 = INput[15];
assign pp_s0_col8_row1 = INput[22];
assign pp_s0_col8_row2 = INput[29];
assign pp_s0_col8_row3 = INput[36];
assign pp_s0_col8_row4 = INput[43];
assign pp_s0_col8_row5 = INput[50];
assign pp_s0_col8_row6 = INput[57];
assign pp_s0_col9_row0 = INput[23];
assign pp_s0_col9_row1 = INput[30];
assign pp_s0_col9_row2 = INput[37];
assign pp_s0_col9_row3 = INput[44];
assign pp_s0_col9_row4 = INput[51];
assign pp_s0_col9_row5 = INput[58];
assign pp_s0_col10_row0 = INput[31];
assign pp_s0_col10_row1 = INput[38];
assign pp_s0_col10_row2 = INput[45];
assign pp_s0_col10_row3 = INput[52];
assign pp_s0_col10_row4 = INput[59];
assign pp_s0_col11_row0 = INput[39];
assign pp_s0_col11_row1 = INput[46];
assign pp_s0_col11_row2 = INput[53];
assign pp_s0_col11_row3 = INput[60];
assign pp_s0_col12_row0 = INput[47];
assign pp_s0_col12_row1 = INput[54];
assign pp_s0_col12_row2 = INput[61];
assign pp_s0_col13_row0 = INput[55];
assign pp_s0_col13_row1 = INput[62];
assign pp_s0_col14_row0 = INput[63];



wire pp_s1_col0_row0;
wire pp_s1_col1_row0;
wire pp_s1_col1_row1;
wire pp_s1_col2_row0;
wire pp_s1_col3_row0;
wire pp_s1_col3_row1;
wire pp_s1_col3_row2;
wire pp_s1_col4_row0;
wire pp_s1_col4_row1;
wire pp_s1_col4_row2;
wire pp_s1_col4_row3;
wire pp_s1_col5_row0;
wire pp_s1_col5_row1;
wire pp_s1_col5_row2;
wire pp_s1_col6_row0;
wire pp_s1_col6_row1;
wire pp_s1_col6_row2;
wire pp_s1_col6_row3;
wire pp_s1_col6_row4;
wire pp_s1_col7_row0;
wire pp_s1_col7_row1;
wire pp_s1_col7_row2;
wire pp_s1_col7_row3;
wire pp_s1_col7_row4;
wire pp_s1_col7_row5;
wire pp_s1_col8_row0;
wire pp_s1_col8_row1;
wire pp_s1_col8_row2;
wire pp_s1_col8_row3;
wire pp_s1_col8_row4;
wire pp_s1_col9_row0;
wire pp_s1_col9_row1;
wire pp_s1_col9_row2;
wire pp_s1_col9_row3;
wire pp_s1_col10_row0;
wire pp_s1_col10_row1;
wire pp_s1_col10_row2;
wire pp_s1_col10_row3;
wire pp_s1_col10_row4;
wire pp_s1_col11_row0;
wire pp_s1_col11_row1;
wire pp_s1_col11_row2;
wire pp_s1_col12_row0;
wire pp_s1_col12_row1;
wire pp_s1_col13_row0;
wire pp_s1_col13_row1;
wire pp_s1_col13_row2;
wire pp_s1_col14_row0;

assign pp_s1_col0_row0 = pp_s0_col0_row0;
assign pp_s1_col1_row0 = pp_s0_col1_row0;
assign pp_s1_col1_row1 = pp_s0_col1_row1;
FullAdder fa_inst_s0_u0 ( .A(pp_s0_col2_row0), .B(pp_s0_col2_row1), .Cin(pp_s0_col2_row2), .Sum(pp_s1_col2_row0), .Cout(pp_s1_col3_row0));
FullAdder fa_inst_s0_u1 ( .A(pp_s0_col3_row0), .B(pp_s0_col3_row1), .Cin(pp_s0_col3_row2), .Sum(pp_s1_col3_row1), .Cout(pp_s1_col4_row0));
assign pp_s1_col3_row2 = pp_s0_col3_row3;
FullAdder fa_inst_s0_u2 ( .A(pp_s0_col4_row0), .B(pp_s0_col4_row1), .Cin(pp_s0_col4_row2), .Sum(pp_s1_col4_row1), .Cout(pp_s1_col5_row0));
assign pp_s1_col4_row2 = pp_s0_col4_row3;
assign pp_s1_col4_row3 = pp_s0_col4_row4;
FullAdder fa_inst_s0_u3 ( .A(pp_s0_col5_row0), .B(pp_s0_col5_row1), .Cin(pp_s0_col5_row2), .Sum(pp_s1_col5_row1), .Cout(pp_s1_col6_row0));
FullAdder fa_inst_s0_u4 ( .A(pp_s0_col5_row3), .B(pp_s0_col5_row4), .Cin(pp_s0_col5_row5), .Sum(pp_s1_col5_row2), .Cout(pp_s1_col6_row1));
FullAdder fa_inst_s0_u5 ( .A(pp_s0_col6_row0), .B(pp_s0_col6_row1), .Cin(pp_s0_col6_row2), .Sum(pp_s1_col6_row2), .Cout(pp_s1_col7_row0));
FullAdder fa_inst_s0_u6 ( .A(pp_s0_col6_row3), .B(pp_s0_col6_row4), .Cin(pp_s0_col6_row5), .Sum(pp_s1_col6_row3), .Cout(pp_s1_col7_row1));
assign pp_s1_col6_row4 = pp_s0_col6_row6;
FullAdder fa_inst_s0_u7 ( .A(pp_s0_col7_row0), .B(pp_s0_col7_row1), .Cin(pp_s0_col7_row2), .Sum(pp_s1_col7_row2), .Cout(pp_s1_col8_row0));
FullAdder fa_inst_s0_u8 ( .A(pp_s0_col7_row3), .B(pp_s0_col7_row4), .Cin(pp_s0_col7_row5), .Sum(pp_s1_col7_row3), .Cout(pp_s1_col8_row1));
assign pp_s1_col7_row4 = pp_s0_col7_row6;
assign pp_s1_col7_row5 = pp_s0_col7_row7;
FullAdder fa_inst_s0_u9 ( .A(pp_s0_col8_row0), .B(pp_s0_col8_row1), .Cin(pp_s0_col8_row2), .Sum(pp_s1_col8_row2), .Cout(pp_s1_col9_row0));
FullAdder fa_inst_s0_u10 ( .A(pp_s0_col8_row3), .B(pp_s0_col8_row4), .Cin(pp_s0_col8_row5), .Sum(pp_s1_col8_row3), .Cout(pp_s1_col9_row1));
assign pp_s1_col8_row4 = pp_s0_col8_row6;
FullAdder fa_inst_s0_u11 ( .A(pp_s0_col9_row0), .B(pp_s0_col9_row1), .Cin(pp_s0_col9_row2), .Sum(pp_s1_col9_row2), .Cout(pp_s1_col10_row0));
FullAdder fa_inst_s0_u12 ( .A(pp_s0_col9_row3), .B(pp_s0_col9_row4), .Cin(pp_s0_col9_row5), .Sum(pp_s1_col9_row3), .Cout(pp_s1_col10_row1));
FullAdder fa_inst_s0_u13 ( .A(pp_s0_col10_row0), .B(pp_s0_col10_row1), .Cin(pp_s0_col10_row2), .Sum(pp_s1_col10_row2), .Cout(pp_s1_col11_row0));
assign pp_s1_col10_row3 = pp_s0_col10_row3;
assign pp_s1_col10_row4 = pp_s0_col10_row4;
FullAdder fa_inst_s0_u14 ( .A(pp_s0_col11_row0), .B(pp_s0_col11_row1), .Cin(pp_s0_col11_row2), .Sum(pp_s1_col11_row1), .Cout(pp_s1_col12_row0));
assign pp_s1_col11_row2 = pp_s0_col11_row3;
FullAdder fa_inst_s0_u15 ( .A(pp_s0_col12_row0), .B(pp_s0_col12_row1), .Cin(pp_s0_col12_row2), .Sum(pp_s1_col12_row1), .Cout(pp_s1_col13_row0));
assign pp_s1_col13_row1 = pp_s0_col13_row0;
assign pp_s1_col13_row2 = pp_s0_col13_row1;
assign pp_s1_col14_row0 = pp_s0_col14_row0;


wire pp_s2_col0_row0;
wire pp_s2_col1_row0;
wire pp_s2_col1_row1;
wire pp_s2_col2_row0;
wire pp_s2_col3_row0;
wire pp_s2_col4_row0;
wire pp_s2_col4_row1;
wire pp_s2_col4_row2;
wire pp_s2_col5_row0;
wire pp_s2_col5_row1;
wire pp_s2_col6_row0;
wire pp_s2_col6_row1;
wire pp_s2_col6_row2;
wire pp_s2_col6_row3;
wire pp_s2_col7_row0;
wire pp_s2_col7_row1;
wire pp_s2_col7_row2;
wire pp_s2_col8_row0;
wire pp_s2_col8_row1;
wire pp_s2_col8_row2;
wire pp_s2_col8_row3;
wire pp_s2_col8_row4;
wire pp_s2_col9_row0;
wire pp_s2_col9_row1;
wire pp_s2_col9_row2;
wire pp_s2_col10_row0;
wire pp_s2_col10_row1;
wire pp_s2_col10_row2;
wire pp_s2_col10_row3;
wire pp_s2_col11_row0;
wire pp_s2_col11_row1;
wire pp_s2_col12_row0;
wire pp_s2_col12_row1;
wire pp_s2_col12_row2;
wire pp_s2_col13_row0;
wire pp_s2_col14_row0;
wire pp_s2_col14_row1;

assign pp_s2_col0_row0 = pp_s1_col0_row0;
assign pp_s2_col1_row0 = pp_s1_col1_row0;
assign pp_s2_col1_row1 = pp_s1_col1_row1;
assign pp_s2_col2_row0 = pp_s1_col2_row0;
FullAdder fa_inst_s1_u0 ( .A(pp_s1_col3_row0), .B(pp_s1_col3_row1), .Cin(pp_s1_col3_row2), .Sum(pp_s2_col3_row0), .Cout(pp_s2_col4_row0));
FullAdder fa_inst_s1_u1 ( .A(pp_s1_col4_row0), .B(pp_s1_col4_row1), .Cin(pp_s1_col4_row2), .Sum(pp_s2_col4_row1), .Cout(pp_s2_col5_row0));
assign pp_s2_col4_row2 = pp_s1_col4_row3;
FullAdder fa_inst_s1_u2 ( .A(pp_s1_col5_row0), .B(pp_s1_col5_row1), .Cin(pp_s1_col5_row2), .Sum(pp_s2_col5_row1), .Cout(pp_s2_col6_row0));
FullAdder fa_inst_s1_u3 ( .A(pp_s1_col6_row0), .B(pp_s1_col6_row1), .Cin(pp_s1_col6_row2), .Sum(pp_s2_col6_row1), .Cout(pp_s2_col7_row0));
assign pp_s2_col6_row2 = pp_s1_col6_row3;
assign pp_s2_col6_row3 = pp_s1_col6_row4;
FullAdder fa_inst_s1_u4 ( .A(pp_s1_col7_row0), .B(pp_s1_col7_row1), .Cin(pp_s1_col7_row2), .Sum(pp_s2_col7_row1), .Cout(pp_s2_col8_row0));
FullAdder fa_inst_s1_u5 ( .A(pp_s1_col7_row3), .B(pp_s1_col7_row4), .Cin(pp_s1_col7_row5), .Sum(pp_s2_col7_row2), .Cout(pp_s2_col8_row1));
FullAdder fa_inst_s1_u6 ( .A(pp_s1_col8_row0), .B(pp_s1_col8_row1), .Cin(pp_s1_col8_row2), .Sum(pp_s2_col8_row2), .Cout(pp_s2_col9_row0));
assign pp_s2_col8_row3 = pp_s1_col8_row3;
assign pp_s2_col8_row4 = pp_s1_col8_row4;
FullAdder fa_inst_s1_u7 ( .A(pp_s1_col9_row0), .B(pp_s1_col9_row1), .Cin(pp_s1_col9_row2), .Sum(pp_s2_col9_row1), .Cout(pp_s2_col10_row0));
assign pp_s2_col9_row2 = pp_s1_col9_row3;
FullAdder fa_inst_s1_u8 ( .A(pp_s1_col10_row0), .B(pp_s1_col10_row1), .Cin(pp_s1_col10_row2), .Sum(pp_s2_col10_row1), .Cout(pp_s2_col11_row0));
assign pp_s2_col10_row2 = pp_s1_col10_row3;
assign pp_s2_col10_row3 = pp_s1_col10_row4;
FullAdder fa_inst_s1_u9 ( .A(pp_s1_col11_row0), .B(pp_s1_col11_row1), .Cin(pp_s1_col11_row2), .Sum(pp_s2_col11_row1), .Cout(pp_s2_col12_row0));
assign pp_s2_col12_row1 = pp_s1_col12_row0;
assign pp_s2_col12_row2 = pp_s1_col12_row1;
FullAdder fa_inst_s1_u10 ( .A(pp_s1_col13_row0), .B(pp_s1_col13_row1), .Cin(pp_s1_col13_row2), .Sum(pp_s2_col13_row0), .Cout(pp_s2_col14_row0));
assign pp_s2_col14_row1 = pp_s1_col14_row0;


wire pp_s3_col0_row0;
wire pp_s3_col1_row0;
wire pp_s3_col1_row1;
wire pp_s3_col2_row0;
wire pp_s3_col3_row0;
wire pp_s3_col4_row0;
wire pp_s3_col5_row0;
wire pp_s3_col5_row1;
wire pp_s3_col5_row2;
wire pp_s3_col6_row0;
wire pp_s3_col6_row1;
wire pp_s3_col7_row0;
wire pp_s3_col7_row1;
wire pp_s3_col8_row0;
wire pp_s3_col8_row1;
wire pp_s3_col8_row2;
wire pp_s3_col8_row3;
wire pp_s3_col9_row0;
wire pp_s3_col9_row1;
wire pp_s3_col10_row0;
wire pp_s3_col10_row1;
wire pp_s3_col10_row2;
wire pp_s3_col11_row0;
wire pp_s3_col11_row1;
wire pp_s3_col11_row2;
wire pp_s3_col12_row0;
wire pp_s3_col13_row0;
wire pp_s3_col13_row1;
wire pp_s3_col14_row0;
wire pp_s3_col14_row1;

assign pp_s3_col0_row0 = pp_s2_col0_row0;
assign pp_s3_col1_row0 = pp_s2_col1_row0;
assign pp_s3_col1_row1 = pp_s2_col1_row1;
assign pp_s3_col2_row0 = pp_s2_col2_row0;
assign pp_s3_col3_row0 = pp_s2_col3_row0;
FullAdder fa_inst_s2_u0 ( .A(pp_s2_col4_row0), .B(pp_s2_col4_row1), .Cin(pp_s2_col4_row2), .Sum(pp_s3_col4_row0), .Cout(pp_s3_col5_row0));
assign pp_s3_col5_row1 = pp_s2_col5_row0;
assign pp_s3_col5_row2 = pp_s2_col5_row1;
FullAdder fa_inst_s2_u1 ( .A(pp_s2_col6_row0), .B(pp_s2_col6_row1), .Cin(pp_s2_col6_row2), .Sum(pp_s3_col6_row0), .Cout(pp_s3_col7_row0));
assign pp_s3_col6_row1 = pp_s2_col6_row3;
FullAdder fa_inst_s2_u2 ( .A(pp_s2_col7_row0), .B(pp_s2_col7_row1), .Cin(pp_s2_col7_row2), .Sum(pp_s3_col7_row1), .Cout(pp_s3_col8_row0));
FullAdder fa_inst_s2_u3 ( .A(pp_s2_col8_row0), .B(pp_s2_col8_row1), .Cin(pp_s2_col8_row2), .Sum(pp_s3_col8_row1), .Cout(pp_s3_col9_row0));
assign pp_s3_col8_row2 = pp_s2_col8_row3;
assign pp_s3_col8_row3 = pp_s2_col8_row4;
FullAdder fa_inst_s2_u4 ( .A(pp_s2_col9_row0), .B(pp_s2_col9_row1), .Cin(pp_s2_col9_row2), .Sum(pp_s3_col9_row1), .Cout(pp_s3_col10_row0));
FullAdder fa_inst_s2_u5 ( .A(pp_s2_col10_row0), .B(pp_s2_col10_row1), .Cin(pp_s2_col10_row2), .Sum(pp_s3_col10_row1), .Cout(pp_s3_col11_row0));
assign pp_s3_col10_row2 = pp_s2_col10_row3;
assign pp_s3_col11_row1 = pp_s2_col11_row0;
assign pp_s3_col11_row2 = pp_s2_col11_row1;
FullAdder fa_inst_s2_u6 ( .A(pp_s2_col12_row0), .B(pp_s2_col12_row1), .Cin(pp_s2_col12_row2), .Sum(pp_s3_col12_row0), .Cout(pp_s3_col13_row0));
assign pp_s3_col13_row1 = pp_s2_col13_row0;
assign pp_s3_col14_row0 = pp_s2_col14_row0;
assign pp_s3_col14_row1 = pp_s2_col14_row1;


wire pp_s4_col0_row0;
wire pp_s4_col1_row0;
wire pp_s4_col1_row1;
wire pp_s4_col2_row0;
wire pp_s4_col3_row0;
wire pp_s4_col4_row0;
wire pp_s4_col5_row0;
wire pp_s4_col6_row0;
wire pp_s4_col6_row1;
wire pp_s4_col6_row2;
wire pp_s4_col7_row0;
wire pp_s4_col7_row1;
wire pp_s4_col8_row0;
wire pp_s4_col8_row1;
wire pp_s4_col9_row0;
wire pp_s4_col9_row1;
wire pp_s4_col9_row2;
wire pp_s4_col10_row0;
wire pp_s4_col11_row0;
wire pp_s4_col11_row1;
wire pp_s4_col12_row0;
wire pp_s4_col12_row1;
wire pp_s4_col13_row0;
wire pp_s4_col13_row1;
wire pp_s4_col14_row0;
wire pp_s4_col14_row1;

assign pp_s4_col0_row0 = pp_s3_col0_row0;
assign pp_s4_col1_row0 = pp_s3_col1_row0;
assign pp_s4_col1_row1 = pp_s3_col1_row1;
assign pp_s4_col2_row0 = pp_s3_col2_row0;
assign pp_s4_col3_row0 = pp_s3_col3_row0;
assign pp_s4_col4_row0 = pp_s3_col4_row0;
FullAdder fa_inst_s3_u0 ( .A(pp_s3_col5_row0), .B(pp_s3_col5_row1), .Cin(pp_s3_col5_row2), .Sum(pp_s4_col5_row0), .Cout(pp_s4_col6_row0));
assign pp_s4_col6_row1 = pp_s3_col6_row0;
assign pp_s4_col6_row2 = pp_s3_col6_row1;
assign pp_s4_col7_row0 = pp_s3_col7_row0;
assign pp_s4_col7_row1 = pp_s3_col7_row1;
FullAdder fa_inst_s3_u1 ( .A(pp_s3_col8_row0), .B(pp_s3_col8_row1), .Cin(pp_s3_col8_row2), .Sum(pp_s4_col8_row0), .Cout(pp_s4_col9_row0));
assign pp_s4_col8_row1 = pp_s3_col8_row3;
assign pp_s4_col9_row1 = pp_s3_col9_row0;
assign pp_s4_col9_row2 = pp_s3_col9_row1;
FullAdder fa_inst_s3_u2 ( .A(pp_s3_col10_row0), .B(pp_s3_col10_row1), .Cin(pp_s3_col10_row2), .Sum(pp_s4_col10_row0), .Cout(pp_s4_col11_row0));
FullAdder fa_inst_s3_u3 ( .A(pp_s3_col11_row0), .B(pp_s3_col11_row1), .Cin(pp_s3_col11_row2), .Sum(pp_s4_col11_row1), .Cout(pp_s4_col12_row0));
assign pp_s4_col12_row1 = pp_s3_col12_row0;
assign pp_s4_col13_row0 = pp_s3_col13_row0;
assign pp_s4_col13_row1 = pp_s3_col13_row1;
assign pp_s4_col14_row0 = pp_s3_col14_row0;
assign pp_s4_col14_row1 = pp_s3_col14_row1;


wire pp_s5_col0_row0;
wire pp_s5_col1_row0;
wire pp_s5_col1_row1;
wire pp_s5_col2_row0;
wire pp_s5_col3_row0;
wire pp_s5_col4_row0;
wire pp_s5_col5_row0;
wire pp_s5_col6_row0;
wire pp_s5_col7_row0;
wire pp_s5_col7_row1;
wire pp_s5_col7_row2;
wire pp_s5_col8_row0;
wire pp_s5_col8_row1;
wire pp_s5_col9_row0;
wire pp_s5_col10_row0;
wire pp_s5_col10_row1;
wire pp_s5_col11_row0;
wire pp_s5_col11_row1;
wire pp_s5_col12_row0;
wire pp_s5_col12_row1;
wire pp_s5_col13_row0;
wire pp_s5_col13_row1;
wire pp_s5_col14_row0;
wire pp_s5_col14_row1;

assign pp_s5_col0_row0 = pp_s4_col0_row0;
assign pp_s5_col1_row0 = pp_s4_col1_row0;
assign pp_s5_col1_row1 = pp_s4_col1_row1;
assign pp_s5_col2_row0 = pp_s4_col2_row0;
assign pp_s5_col3_row0 = pp_s4_col3_row0;
assign pp_s5_col4_row0 = pp_s4_col4_row0;
assign pp_s5_col5_row0 = pp_s4_col5_row0;
FullAdder fa_inst_s4_u0 ( .A(pp_s4_col6_row0), .B(pp_s4_col6_row1), .Cin(pp_s4_col6_row2), .Sum(pp_s5_col6_row0), .Cout(pp_s5_col7_row0));
assign pp_s5_col7_row1 = pp_s4_col7_row0;
assign pp_s5_col7_row2 = pp_s4_col7_row1;
assign pp_s5_col8_row0 = pp_s4_col8_row0;
assign pp_s5_col8_row1 = pp_s4_col8_row1;
FullAdder fa_inst_s4_u1 ( .A(pp_s4_col9_row0), .B(pp_s4_col9_row1), .Cin(pp_s4_col9_row2), .Sum(pp_s5_col9_row0), .Cout(pp_s5_col10_row0));
assign pp_s5_col10_row1 = pp_s4_col10_row0;
assign pp_s5_col11_row0 = pp_s4_col11_row0;
assign pp_s5_col11_row1 = pp_s4_col11_row1;
assign pp_s5_col12_row0 = pp_s4_col12_row0;
assign pp_s5_col12_row1 = pp_s4_col12_row1;
assign pp_s5_col13_row0 = pp_s4_col13_row0;
assign pp_s5_col13_row1 = pp_s4_col13_row1;
assign pp_s5_col14_row0 = pp_s4_col14_row0;
assign pp_s5_col14_row1 = pp_s4_col14_row1;


wire pp_s6_col0_row0;
wire pp_s6_col1_row0;
wire pp_s6_col1_row1;
wire pp_s6_col2_row0;
wire pp_s6_col3_row0;
wire pp_s6_col4_row0;
wire pp_s6_col5_row0;
wire pp_s6_col6_row0;
wire pp_s6_col7_row0;
wire pp_s6_col8_row0;
wire pp_s6_col8_row1;
wire pp_s6_col8_row2;
wire pp_s6_col9_row0;
wire pp_s6_col10_row0;
wire pp_s6_col10_row1;
wire pp_s6_col11_row0;
wire pp_s6_col11_row1;
wire pp_s6_col12_row0;
wire pp_s6_col12_row1;
wire pp_s6_col13_row0;
wire pp_s6_col13_row1;
wire pp_s6_col14_row0;
wire pp_s6_col14_row1;

assign pp_s6_col0_row0 = pp_s5_col0_row0;
assign pp_s6_col1_row0 = pp_s5_col1_row0;
assign pp_s6_col1_row1 = pp_s5_col1_row1;
assign pp_s6_col2_row0 = pp_s5_col2_row0;
assign pp_s6_col3_row0 = pp_s5_col3_row0;
assign pp_s6_col4_row0 = pp_s5_col4_row0;
assign pp_s6_col5_row0 = pp_s5_col5_row0;
assign pp_s6_col6_row0 = pp_s5_col6_row0;
FullAdder fa_inst_s5_u0 ( .A(pp_s5_col7_row0), .B(pp_s5_col7_row1), .Cin(pp_s5_col7_row2), .Sum(pp_s6_col7_row0), .Cout(pp_s6_col8_row0));
assign pp_s6_col8_row1 = pp_s5_col8_row0;
assign pp_s6_col8_row2 = pp_s5_col8_row1;
assign pp_s6_col9_row0 = pp_s5_col9_row0;
assign pp_s6_col10_row0 = pp_s5_col10_row0;
assign pp_s6_col10_row1 = pp_s5_col10_row1;
assign pp_s6_col11_row0 = pp_s5_col11_row0;
assign pp_s6_col11_row1 = pp_s5_col11_row1;
assign pp_s6_col12_row0 = pp_s5_col12_row0;
assign pp_s6_col12_row1 = pp_s5_col12_row1;
assign pp_s6_col13_row0 = pp_s5_col13_row0;
assign pp_s6_col13_row1 = pp_s5_col13_row1;
assign pp_s6_col14_row0 = pp_s5_col14_row0;
assign pp_s6_col14_row1 = pp_s5_col14_row1;


wire pp_s7_col0_row0;
wire pp_s7_col1_row0;
wire pp_s7_col1_row1;
wire pp_s7_col2_row0;
wire pp_s7_col3_row0;
wire pp_s7_col4_row0;
wire pp_s7_col5_row0;
wire pp_s7_col6_row0;
wire pp_s7_col7_row0;
wire pp_s7_col8_row0;
wire pp_s7_col9_row0;
wire pp_s7_col9_row1;
wire pp_s7_col10_row0;
wire pp_s7_col10_row1;
wire pp_s7_col11_row0;
wire pp_s7_col11_row1;
wire pp_s7_col12_row0;
wire pp_s7_col12_row1;
wire pp_s7_col13_row0;
wire pp_s7_col13_row1;
wire pp_s7_col14_row0;
wire pp_s7_col14_row1;

assign pp_s7_col0_row0 = pp_s6_col0_row0;
assign pp_s7_col1_row0 = pp_s6_col1_row0;
assign pp_s7_col1_row1 = pp_s6_col1_row1;
assign pp_s7_col2_row0 = pp_s6_col2_row0;
assign pp_s7_col3_row0 = pp_s6_col3_row0;
assign pp_s7_col4_row0 = pp_s6_col4_row0;
assign pp_s7_col5_row0 = pp_s6_col5_row0;
assign pp_s7_col6_row0 = pp_s6_col6_row0;
assign pp_s7_col7_row0 = pp_s6_col7_row0;
FullAdder fa_inst_s6_u0 ( .A(pp_s6_col8_row0), .B(pp_s6_col8_row1), .Cin(pp_s6_col8_row2), .Sum(pp_s7_col8_row0), .Cout(pp_s7_col9_row0));
assign pp_s7_col9_row1 = pp_s6_col9_row0;
assign pp_s7_col10_row0 = pp_s6_col10_row0;
assign pp_s7_col10_row1 = pp_s6_col10_row1;
assign pp_s7_col11_row0 = pp_s6_col11_row0;
assign pp_s7_col11_row1 = pp_s6_col11_row1;
assign pp_s7_col12_row0 = pp_s6_col12_row0;
assign pp_s7_col12_row1 = pp_s6_col12_row1;
assign pp_s7_col13_row0 = pp_s6_col13_row0;
assign pp_s7_col13_row1 = pp_s6_col13_row1;
assign pp_s7_col14_row0 = pp_s6_col14_row0;
assign pp_s7_col14_row1 = pp_s6_col14_row1;

assign WALLACEout[0][0] = pp_s7_col0_row0;
assign WALLACEout[0][1] = pp_s7_col1_row0;
assign WALLACEout[1][1] = pp_s7_col1_row1;
assign WALLACEout[0][2] = pp_s7_col2_row0;
assign WALLACEout[0][3] = pp_s7_col3_row0;
assign WALLACEout[0][4] = pp_s7_col4_row0;
assign WALLACEout[0][5] = pp_s7_col5_row0;
assign WALLACEout[0][6] = pp_s7_col6_row0;
assign WALLACEout[0][7] = pp_s7_col7_row0;
assign WALLACEout[0][8] = pp_s7_col8_row0;
assign WALLACEout[0][9] = pp_s7_col9_row0;
assign WALLACEout[1][9] = pp_s7_col9_row1;
assign WALLACEout[0][10] = pp_s7_col10_row0;
assign WALLACEout[1][10] = pp_s7_col10_row1;
assign WALLACEout[0][11] = pp_s7_col11_row0;
assign WALLACEout[1][11] = pp_s7_col11_row1;
assign WALLACEout[0][12] = pp_s7_col12_row0;
assign WALLACEout[1][12] = pp_s7_col12_row1;
assign WALLACEout[0][13] = pp_s7_col13_row0;
assign WALLACEout[1][13] = pp_s7_col13_row1;
assign WALLACEout[0][14] = pp_s7_col14_row0;
assign WALLACEout[1][14] = pp_s7_col14_row1;

endmodule;
